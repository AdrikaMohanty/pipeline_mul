magic
tech sky130A
magscale 1 2
timestamp 1700931726
<< obsli1 >>
rect 1104 2159 318872 317713
<< obsm1 >>
rect 1104 2128 318872 317744
<< metal2 >>
rect 5354 319200 5410 320000
rect 14186 319200 14242 320000
rect 23018 319200 23074 320000
rect 31850 319200 31906 320000
rect 40682 319200 40738 320000
rect 49514 319200 49570 320000
rect 58346 319200 58402 320000
rect 67178 319200 67234 320000
rect 76010 319200 76066 320000
rect 84842 319200 84898 320000
rect 93674 319200 93730 320000
rect 102506 319200 102562 320000
rect 111338 319200 111394 320000
rect 120170 319200 120226 320000
rect 129002 319200 129058 320000
rect 137834 319200 137890 320000
rect 146666 319200 146722 320000
rect 155498 319200 155554 320000
rect 164330 319200 164386 320000
rect 173162 319200 173218 320000
rect 181994 319200 182050 320000
rect 190826 319200 190882 320000
rect 199658 319200 199714 320000
rect 208490 319200 208546 320000
rect 217322 319200 217378 320000
rect 226154 319200 226210 320000
rect 234986 319200 235042 320000
rect 243818 319200 243874 320000
rect 252650 319200 252706 320000
rect 261482 319200 261538 320000
rect 270314 319200 270370 320000
rect 279146 319200 279202 320000
rect 287978 319200 288034 320000
rect 296810 319200 296866 320000
rect 305642 319200 305698 320000
rect 314474 319200 314530 320000
rect 1214 0 1270 800
rect 1858 0 1914 800
rect 2502 0 2558 800
rect 3146 0 3202 800
rect 3790 0 3846 800
rect 4434 0 4490 800
rect 5078 0 5134 800
rect 5722 0 5778 800
rect 6366 0 6422 800
rect 7010 0 7066 800
rect 7654 0 7710 800
rect 8298 0 8354 800
rect 8942 0 8998 800
rect 9586 0 9642 800
rect 10230 0 10286 800
rect 10874 0 10930 800
rect 11518 0 11574 800
rect 12162 0 12218 800
rect 12806 0 12862 800
rect 13450 0 13506 800
rect 14094 0 14150 800
rect 14738 0 14794 800
rect 15382 0 15438 800
rect 16026 0 16082 800
rect 16670 0 16726 800
rect 17314 0 17370 800
rect 17958 0 18014 800
rect 18602 0 18658 800
rect 19246 0 19302 800
rect 19890 0 19946 800
rect 20534 0 20590 800
rect 21178 0 21234 800
rect 21822 0 21878 800
rect 22466 0 22522 800
rect 23110 0 23166 800
rect 23754 0 23810 800
rect 24398 0 24454 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 26974 0 27030 800
rect 27618 0 27674 800
rect 28262 0 28318 800
rect 28906 0 28962 800
rect 29550 0 29606 800
rect 30194 0 30250 800
rect 30838 0 30894 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33414 0 33470 800
rect 34058 0 34114 800
rect 34702 0 34758 800
rect 35346 0 35402 800
rect 35990 0 36046 800
rect 36634 0 36690 800
rect 37278 0 37334 800
rect 37922 0 37978 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39854 0 39910 800
rect 40498 0 40554 800
rect 41142 0 41198 800
rect 41786 0 41842 800
rect 42430 0 42486 800
rect 43074 0 43130 800
rect 43718 0 43774 800
rect 44362 0 44418 800
rect 45006 0 45062 800
rect 45650 0 45706 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47582 0 47638 800
rect 48226 0 48282 800
rect 48870 0 48926 800
rect 49514 0 49570 800
rect 50158 0 50214 800
rect 50802 0 50858 800
rect 51446 0 51502 800
rect 52090 0 52146 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 54022 0 54078 800
rect 54666 0 54722 800
rect 55310 0 55366 800
rect 55954 0 56010 800
rect 56598 0 56654 800
rect 57242 0 57298 800
rect 57886 0 57942 800
rect 58530 0 58586 800
rect 59174 0 59230 800
rect 59818 0 59874 800
rect 60462 0 60518 800
rect 61106 0 61162 800
rect 61750 0 61806 800
rect 62394 0 62450 800
rect 63038 0 63094 800
rect 63682 0 63738 800
rect 64326 0 64382 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66258 0 66314 800
rect 66902 0 66958 800
rect 67546 0 67602 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69478 0 69534 800
rect 70122 0 70178 800
rect 70766 0 70822 800
rect 71410 0 71466 800
rect 72054 0 72110 800
rect 72698 0 72754 800
rect 73342 0 73398 800
rect 73986 0 74042 800
rect 74630 0 74686 800
rect 75274 0 75330 800
rect 75918 0 75974 800
rect 76562 0 76618 800
rect 77206 0 77262 800
rect 77850 0 77906 800
rect 78494 0 78550 800
rect 79138 0 79194 800
rect 79782 0 79838 800
rect 80426 0 80482 800
rect 81070 0 81126 800
rect 81714 0 81770 800
rect 82358 0 82414 800
rect 83002 0 83058 800
rect 83646 0 83702 800
rect 84290 0 84346 800
rect 84934 0 84990 800
rect 85578 0 85634 800
rect 86222 0 86278 800
rect 86866 0 86922 800
rect 87510 0 87566 800
rect 88154 0 88210 800
rect 88798 0 88854 800
rect 89442 0 89498 800
rect 90086 0 90142 800
rect 90730 0 90786 800
rect 91374 0 91430 800
rect 92018 0 92074 800
rect 92662 0 92718 800
rect 93306 0 93362 800
rect 93950 0 94006 800
rect 94594 0 94650 800
rect 95238 0 95294 800
rect 95882 0 95938 800
rect 96526 0 96582 800
rect 97170 0 97226 800
rect 97814 0 97870 800
rect 98458 0 98514 800
rect 99102 0 99158 800
rect 99746 0 99802 800
rect 100390 0 100446 800
rect 101034 0 101090 800
rect 101678 0 101734 800
rect 102322 0 102378 800
rect 102966 0 103022 800
rect 103610 0 103666 800
rect 104254 0 104310 800
rect 104898 0 104954 800
rect 105542 0 105598 800
rect 106186 0 106242 800
rect 106830 0 106886 800
rect 107474 0 107530 800
rect 108118 0 108174 800
rect 108762 0 108818 800
rect 109406 0 109462 800
rect 110050 0 110106 800
rect 110694 0 110750 800
rect 111338 0 111394 800
rect 111982 0 112038 800
rect 112626 0 112682 800
rect 113270 0 113326 800
rect 113914 0 113970 800
rect 114558 0 114614 800
rect 115202 0 115258 800
rect 115846 0 115902 800
rect 116490 0 116546 800
rect 117134 0 117190 800
rect 117778 0 117834 800
rect 118422 0 118478 800
rect 119066 0 119122 800
rect 119710 0 119766 800
rect 120354 0 120410 800
rect 120998 0 121054 800
rect 121642 0 121698 800
rect 122286 0 122342 800
rect 122930 0 122986 800
rect 123574 0 123630 800
rect 124218 0 124274 800
rect 124862 0 124918 800
rect 125506 0 125562 800
rect 126150 0 126206 800
rect 126794 0 126850 800
rect 127438 0 127494 800
rect 128082 0 128138 800
rect 128726 0 128782 800
rect 129370 0 129426 800
rect 130014 0 130070 800
rect 130658 0 130714 800
rect 131302 0 131358 800
rect 131946 0 132002 800
rect 132590 0 132646 800
rect 133234 0 133290 800
rect 133878 0 133934 800
rect 134522 0 134578 800
rect 135166 0 135222 800
rect 135810 0 135866 800
rect 136454 0 136510 800
rect 137098 0 137154 800
rect 137742 0 137798 800
rect 138386 0 138442 800
rect 139030 0 139086 800
rect 139674 0 139730 800
rect 140318 0 140374 800
rect 140962 0 141018 800
rect 141606 0 141662 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143538 0 143594 800
rect 144182 0 144238 800
rect 144826 0 144882 800
rect 145470 0 145526 800
rect 146114 0 146170 800
rect 146758 0 146814 800
rect 147402 0 147458 800
rect 148046 0 148102 800
rect 148690 0 148746 800
rect 149334 0 149390 800
rect 149978 0 150034 800
rect 150622 0 150678 800
rect 151266 0 151322 800
rect 151910 0 151966 800
rect 152554 0 152610 800
rect 153198 0 153254 800
rect 153842 0 153898 800
rect 154486 0 154542 800
rect 155130 0 155186 800
rect 155774 0 155830 800
rect 156418 0 156474 800
rect 157062 0 157118 800
rect 157706 0 157762 800
rect 158350 0 158406 800
rect 158994 0 159050 800
rect 159638 0 159694 800
rect 160282 0 160338 800
rect 160926 0 160982 800
rect 161570 0 161626 800
rect 162214 0 162270 800
rect 162858 0 162914 800
rect 163502 0 163558 800
rect 164146 0 164202 800
rect 164790 0 164846 800
rect 165434 0 165490 800
rect 166078 0 166134 800
rect 166722 0 166778 800
rect 167366 0 167422 800
rect 168010 0 168066 800
rect 168654 0 168710 800
rect 169298 0 169354 800
rect 169942 0 169998 800
rect 170586 0 170642 800
rect 171230 0 171286 800
rect 171874 0 171930 800
rect 172518 0 172574 800
rect 173162 0 173218 800
rect 173806 0 173862 800
rect 174450 0 174506 800
rect 175094 0 175150 800
rect 175738 0 175794 800
rect 176382 0 176438 800
rect 177026 0 177082 800
rect 177670 0 177726 800
rect 178314 0 178370 800
rect 178958 0 179014 800
rect 179602 0 179658 800
rect 180246 0 180302 800
rect 180890 0 180946 800
rect 181534 0 181590 800
rect 182178 0 182234 800
rect 182822 0 182878 800
rect 183466 0 183522 800
rect 184110 0 184166 800
rect 184754 0 184810 800
rect 185398 0 185454 800
rect 186042 0 186098 800
rect 186686 0 186742 800
rect 187330 0 187386 800
rect 187974 0 188030 800
rect 188618 0 188674 800
rect 189262 0 189318 800
rect 189906 0 189962 800
rect 190550 0 190606 800
rect 191194 0 191250 800
rect 191838 0 191894 800
rect 192482 0 192538 800
rect 193126 0 193182 800
rect 193770 0 193826 800
rect 194414 0 194470 800
rect 195058 0 195114 800
rect 195702 0 195758 800
rect 196346 0 196402 800
rect 196990 0 197046 800
rect 197634 0 197690 800
rect 198278 0 198334 800
rect 198922 0 198978 800
rect 199566 0 199622 800
rect 200210 0 200266 800
rect 200854 0 200910 800
rect 201498 0 201554 800
rect 202142 0 202198 800
rect 202786 0 202842 800
rect 203430 0 203486 800
rect 204074 0 204130 800
rect 204718 0 204774 800
rect 205362 0 205418 800
rect 206006 0 206062 800
rect 206650 0 206706 800
rect 207294 0 207350 800
rect 207938 0 207994 800
rect 208582 0 208638 800
rect 209226 0 209282 800
rect 209870 0 209926 800
rect 210514 0 210570 800
rect 211158 0 211214 800
rect 211802 0 211858 800
rect 212446 0 212502 800
rect 213090 0 213146 800
rect 213734 0 213790 800
rect 214378 0 214434 800
rect 215022 0 215078 800
rect 215666 0 215722 800
rect 216310 0 216366 800
rect 216954 0 217010 800
rect 217598 0 217654 800
rect 218242 0 218298 800
rect 218886 0 218942 800
rect 219530 0 219586 800
rect 220174 0 220230 800
rect 220818 0 220874 800
rect 221462 0 221518 800
rect 222106 0 222162 800
rect 222750 0 222806 800
rect 223394 0 223450 800
rect 224038 0 224094 800
rect 224682 0 224738 800
rect 225326 0 225382 800
rect 225970 0 226026 800
rect 226614 0 226670 800
rect 227258 0 227314 800
rect 227902 0 227958 800
rect 228546 0 228602 800
rect 229190 0 229246 800
rect 229834 0 229890 800
rect 230478 0 230534 800
rect 231122 0 231178 800
rect 231766 0 231822 800
rect 232410 0 232466 800
rect 233054 0 233110 800
rect 233698 0 233754 800
rect 234342 0 234398 800
rect 234986 0 235042 800
rect 235630 0 235686 800
rect 236274 0 236330 800
rect 236918 0 236974 800
rect 237562 0 237618 800
rect 238206 0 238262 800
rect 238850 0 238906 800
rect 239494 0 239550 800
rect 240138 0 240194 800
rect 240782 0 240838 800
rect 241426 0 241482 800
rect 242070 0 242126 800
rect 242714 0 242770 800
rect 243358 0 243414 800
rect 244002 0 244058 800
rect 244646 0 244702 800
rect 245290 0 245346 800
rect 245934 0 245990 800
rect 246578 0 246634 800
rect 247222 0 247278 800
rect 247866 0 247922 800
rect 248510 0 248566 800
rect 249154 0 249210 800
rect 249798 0 249854 800
rect 250442 0 250498 800
rect 251086 0 251142 800
rect 251730 0 251786 800
rect 252374 0 252430 800
rect 253018 0 253074 800
rect 253662 0 253718 800
rect 254306 0 254362 800
rect 254950 0 255006 800
rect 255594 0 255650 800
rect 256238 0 256294 800
rect 256882 0 256938 800
rect 257526 0 257582 800
rect 258170 0 258226 800
rect 258814 0 258870 800
rect 259458 0 259514 800
rect 260102 0 260158 800
rect 260746 0 260802 800
rect 261390 0 261446 800
rect 262034 0 262090 800
rect 262678 0 262734 800
rect 263322 0 263378 800
rect 263966 0 264022 800
rect 264610 0 264666 800
rect 265254 0 265310 800
rect 265898 0 265954 800
rect 266542 0 266598 800
rect 267186 0 267242 800
rect 267830 0 267886 800
rect 268474 0 268530 800
rect 269118 0 269174 800
rect 269762 0 269818 800
rect 270406 0 270462 800
rect 271050 0 271106 800
rect 271694 0 271750 800
rect 272338 0 272394 800
rect 272982 0 273038 800
rect 273626 0 273682 800
rect 274270 0 274326 800
rect 274914 0 274970 800
rect 275558 0 275614 800
rect 276202 0 276258 800
rect 276846 0 276902 800
rect 277490 0 277546 800
rect 278134 0 278190 800
rect 278778 0 278834 800
rect 279422 0 279478 800
rect 280066 0 280122 800
rect 280710 0 280766 800
rect 281354 0 281410 800
rect 281998 0 282054 800
rect 282642 0 282698 800
rect 283286 0 283342 800
rect 283930 0 283986 800
rect 284574 0 284630 800
rect 285218 0 285274 800
rect 285862 0 285918 800
rect 286506 0 286562 800
rect 287150 0 287206 800
rect 287794 0 287850 800
rect 288438 0 288494 800
rect 289082 0 289138 800
rect 289726 0 289782 800
rect 290370 0 290426 800
rect 291014 0 291070 800
rect 291658 0 291714 800
rect 292302 0 292358 800
rect 292946 0 293002 800
rect 293590 0 293646 800
rect 294234 0 294290 800
rect 294878 0 294934 800
rect 295522 0 295578 800
rect 296166 0 296222 800
rect 296810 0 296866 800
rect 297454 0 297510 800
rect 298098 0 298154 800
rect 298742 0 298798 800
rect 299386 0 299442 800
rect 300030 0 300086 800
rect 300674 0 300730 800
rect 301318 0 301374 800
rect 301962 0 302018 800
rect 302606 0 302662 800
rect 303250 0 303306 800
rect 303894 0 303950 800
rect 304538 0 304594 800
rect 305182 0 305238 800
rect 305826 0 305882 800
rect 306470 0 306526 800
rect 307114 0 307170 800
rect 307758 0 307814 800
rect 308402 0 308458 800
rect 309046 0 309102 800
rect 309690 0 309746 800
rect 310334 0 310390 800
rect 310978 0 311034 800
rect 311622 0 311678 800
rect 312266 0 312322 800
rect 312910 0 312966 800
rect 313554 0 313610 800
rect 314198 0 314254 800
rect 314842 0 314898 800
rect 315486 0 315542 800
rect 316130 0 316186 800
rect 316774 0 316830 800
rect 317418 0 317474 800
rect 318062 0 318118 800
rect 318706 0 318762 800
<< obsm2 >>
rect 1216 319144 5298 319200
rect 5466 319144 14130 319200
rect 14298 319144 22962 319200
rect 23130 319144 31794 319200
rect 31962 319144 40626 319200
rect 40794 319144 49458 319200
rect 49626 319144 58290 319200
rect 58458 319144 67122 319200
rect 67290 319144 75954 319200
rect 76122 319144 84786 319200
rect 84954 319144 93618 319200
rect 93786 319144 102450 319200
rect 102618 319144 111282 319200
rect 111450 319144 120114 319200
rect 120282 319144 128946 319200
rect 129114 319144 137778 319200
rect 137946 319144 146610 319200
rect 146778 319144 155442 319200
rect 155610 319144 164274 319200
rect 164442 319144 173106 319200
rect 173274 319144 181938 319200
rect 182106 319144 190770 319200
rect 190938 319144 199602 319200
rect 199770 319144 208434 319200
rect 208602 319144 217266 319200
rect 217434 319144 226098 319200
rect 226266 319144 234930 319200
rect 235098 319144 243762 319200
rect 243930 319144 252594 319200
rect 252762 319144 261426 319200
rect 261594 319144 270258 319200
rect 270426 319144 279090 319200
rect 279258 319144 287922 319200
rect 288090 319144 296754 319200
rect 296922 319144 305586 319200
rect 305754 319144 314418 319200
rect 314586 319144 318760 319200
rect 1216 856 318760 319144
rect 1326 734 1802 856
rect 1970 734 2446 856
rect 2614 734 3090 856
rect 3258 734 3734 856
rect 3902 734 4378 856
rect 4546 734 5022 856
rect 5190 734 5666 856
rect 5834 734 6310 856
rect 6478 734 6954 856
rect 7122 734 7598 856
rect 7766 734 8242 856
rect 8410 734 8886 856
rect 9054 734 9530 856
rect 9698 734 10174 856
rect 10342 734 10818 856
rect 10986 734 11462 856
rect 11630 734 12106 856
rect 12274 734 12750 856
rect 12918 734 13394 856
rect 13562 734 14038 856
rect 14206 734 14682 856
rect 14850 734 15326 856
rect 15494 734 15970 856
rect 16138 734 16614 856
rect 16782 734 17258 856
rect 17426 734 17902 856
rect 18070 734 18546 856
rect 18714 734 19190 856
rect 19358 734 19834 856
rect 20002 734 20478 856
rect 20646 734 21122 856
rect 21290 734 21766 856
rect 21934 734 22410 856
rect 22578 734 23054 856
rect 23222 734 23698 856
rect 23866 734 24342 856
rect 24510 734 24986 856
rect 25154 734 25630 856
rect 25798 734 26274 856
rect 26442 734 26918 856
rect 27086 734 27562 856
rect 27730 734 28206 856
rect 28374 734 28850 856
rect 29018 734 29494 856
rect 29662 734 30138 856
rect 30306 734 30782 856
rect 30950 734 31426 856
rect 31594 734 32070 856
rect 32238 734 32714 856
rect 32882 734 33358 856
rect 33526 734 34002 856
rect 34170 734 34646 856
rect 34814 734 35290 856
rect 35458 734 35934 856
rect 36102 734 36578 856
rect 36746 734 37222 856
rect 37390 734 37866 856
rect 38034 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39798 856
rect 39966 734 40442 856
rect 40610 734 41086 856
rect 41254 734 41730 856
rect 41898 734 42374 856
rect 42542 734 43018 856
rect 43186 734 43662 856
rect 43830 734 44306 856
rect 44474 734 44950 856
rect 45118 734 45594 856
rect 45762 734 46238 856
rect 46406 734 46882 856
rect 47050 734 47526 856
rect 47694 734 48170 856
rect 48338 734 48814 856
rect 48982 734 49458 856
rect 49626 734 50102 856
rect 50270 734 50746 856
rect 50914 734 51390 856
rect 51558 734 52034 856
rect 52202 734 52678 856
rect 52846 734 53322 856
rect 53490 734 53966 856
rect 54134 734 54610 856
rect 54778 734 55254 856
rect 55422 734 55898 856
rect 56066 734 56542 856
rect 56710 734 57186 856
rect 57354 734 57830 856
rect 57998 734 58474 856
rect 58642 734 59118 856
rect 59286 734 59762 856
rect 59930 734 60406 856
rect 60574 734 61050 856
rect 61218 734 61694 856
rect 61862 734 62338 856
rect 62506 734 62982 856
rect 63150 734 63626 856
rect 63794 734 64270 856
rect 64438 734 64914 856
rect 65082 734 65558 856
rect 65726 734 66202 856
rect 66370 734 66846 856
rect 67014 734 67490 856
rect 67658 734 68134 856
rect 68302 734 68778 856
rect 68946 734 69422 856
rect 69590 734 70066 856
rect 70234 734 70710 856
rect 70878 734 71354 856
rect 71522 734 71998 856
rect 72166 734 72642 856
rect 72810 734 73286 856
rect 73454 734 73930 856
rect 74098 734 74574 856
rect 74742 734 75218 856
rect 75386 734 75862 856
rect 76030 734 76506 856
rect 76674 734 77150 856
rect 77318 734 77794 856
rect 77962 734 78438 856
rect 78606 734 79082 856
rect 79250 734 79726 856
rect 79894 734 80370 856
rect 80538 734 81014 856
rect 81182 734 81658 856
rect 81826 734 82302 856
rect 82470 734 82946 856
rect 83114 734 83590 856
rect 83758 734 84234 856
rect 84402 734 84878 856
rect 85046 734 85522 856
rect 85690 734 86166 856
rect 86334 734 86810 856
rect 86978 734 87454 856
rect 87622 734 88098 856
rect 88266 734 88742 856
rect 88910 734 89386 856
rect 89554 734 90030 856
rect 90198 734 90674 856
rect 90842 734 91318 856
rect 91486 734 91962 856
rect 92130 734 92606 856
rect 92774 734 93250 856
rect 93418 734 93894 856
rect 94062 734 94538 856
rect 94706 734 95182 856
rect 95350 734 95826 856
rect 95994 734 96470 856
rect 96638 734 97114 856
rect 97282 734 97758 856
rect 97926 734 98402 856
rect 98570 734 99046 856
rect 99214 734 99690 856
rect 99858 734 100334 856
rect 100502 734 100978 856
rect 101146 734 101622 856
rect 101790 734 102266 856
rect 102434 734 102910 856
rect 103078 734 103554 856
rect 103722 734 104198 856
rect 104366 734 104842 856
rect 105010 734 105486 856
rect 105654 734 106130 856
rect 106298 734 106774 856
rect 106942 734 107418 856
rect 107586 734 108062 856
rect 108230 734 108706 856
rect 108874 734 109350 856
rect 109518 734 109994 856
rect 110162 734 110638 856
rect 110806 734 111282 856
rect 111450 734 111926 856
rect 112094 734 112570 856
rect 112738 734 113214 856
rect 113382 734 113858 856
rect 114026 734 114502 856
rect 114670 734 115146 856
rect 115314 734 115790 856
rect 115958 734 116434 856
rect 116602 734 117078 856
rect 117246 734 117722 856
rect 117890 734 118366 856
rect 118534 734 119010 856
rect 119178 734 119654 856
rect 119822 734 120298 856
rect 120466 734 120942 856
rect 121110 734 121586 856
rect 121754 734 122230 856
rect 122398 734 122874 856
rect 123042 734 123518 856
rect 123686 734 124162 856
rect 124330 734 124806 856
rect 124974 734 125450 856
rect 125618 734 126094 856
rect 126262 734 126738 856
rect 126906 734 127382 856
rect 127550 734 128026 856
rect 128194 734 128670 856
rect 128838 734 129314 856
rect 129482 734 129958 856
rect 130126 734 130602 856
rect 130770 734 131246 856
rect 131414 734 131890 856
rect 132058 734 132534 856
rect 132702 734 133178 856
rect 133346 734 133822 856
rect 133990 734 134466 856
rect 134634 734 135110 856
rect 135278 734 135754 856
rect 135922 734 136398 856
rect 136566 734 137042 856
rect 137210 734 137686 856
rect 137854 734 138330 856
rect 138498 734 138974 856
rect 139142 734 139618 856
rect 139786 734 140262 856
rect 140430 734 140906 856
rect 141074 734 141550 856
rect 141718 734 142194 856
rect 142362 734 142838 856
rect 143006 734 143482 856
rect 143650 734 144126 856
rect 144294 734 144770 856
rect 144938 734 145414 856
rect 145582 734 146058 856
rect 146226 734 146702 856
rect 146870 734 147346 856
rect 147514 734 147990 856
rect 148158 734 148634 856
rect 148802 734 149278 856
rect 149446 734 149922 856
rect 150090 734 150566 856
rect 150734 734 151210 856
rect 151378 734 151854 856
rect 152022 734 152498 856
rect 152666 734 153142 856
rect 153310 734 153786 856
rect 153954 734 154430 856
rect 154598 734 155074 856
rect 155242 734 155718 856
rect 155886 734 156362 856
rect 156530 734 157006 856
rect 157174 734 157650 856
rect 157818 734 158294 856
rect 158462 734 158938 856
rect 159106 734 159582 856
rect 159750 734 160226 856
rect 160394 734 160870 856
rect 161038 734 161514 856
rect 161682 734 162158 856
rect 162326 734 162802 856
rect 162970 734 163446 856
rect 163614 734 164090 856
rect 164258 734 164734 856
rect 164902 734 165378 856
rect 165546 734 166022 856
rect 166190 734 166666 856
rect 166834 734 167310 856
rect 167478 734 167954 856
rect 168122 734 168598 856
rect 168766 734 169242 856
rect 169410 734 169886 856
rect 170054 734 170530 856
rect 170698 734 171174 856
rect 171342 734 171818 856
rect 171986 734 172462 856
rect 172630 734 173106 856
rect 173274 734 173750 856
rect 173918 734 174394 856
rect 174562 734 175038 856
rect 175206 734 175682 856
rect 175850 734 176326 856
rect 176494 734 176970 856
rect 177138 734 177614 856
rect 177782 734 178258 856
rect 178426 734 178902 856
rect 179070 734 179546 856
rect 179714 734 180190 856
rect 180358 734 180834 856
rect 181002 734 181478 856
rect 181646 734 182122 856
rect 182290 734 182766 856
rect 182934 734 183410 856
rect 183578 734 184054 856
rect 184222 734 184698 856
rect 184866 734 185342 856
rect 185510 734 185986 856
rect 186154 734 186630 856
rect 186798 734 187274 856
rect 187442 734 187918 856
rect 188086 734 188562 856
rect 188730 734 189206 856
rect 189374 734 189850 856
rect 190018 734 190494 856
rect 190662 734 191138 856
rect 191306 734 191782 856
rect 191950 734 192426 856
rect 192594 734 193070 856
rect 193238 734 193714 856
rect 193882 734 194358 856
rect 194526 734 195002 856
rect 195170 734 195646 856
rect 195814 734 196290 856
rect 196458 734 196934 856
rect 197102 734 197578 856
rect 197746 734 198222 856
rect 198390 734 198866 856
rect 199034 734 199510 856
rect 199678 734 200154 856
rect 200322 734 200798 856
rect 200966 734 201442 856
rect 201610 734 202086 856
rect 202254 734 202730 856
rect 202898 734 203374 856
rect 203542 734 204018 856
rect 204186 734 204662 856
rect 204830 734 205306 856
rect 205474 734 205950 856
rect 206118 734 206594 856
rect 206762 734 207238 856
rect 207406 734 207882 856
rect 208050 734 208526 856
rect 208694 734 209170 856
rect 209338 734 209814 856
rect 209982 734 210458 856
rect 210626 734 211102 856
rect 211270 734 211746 856
rect 211914 734 212390 856
rect 212558 734 213034 856
rect 213202 734 213678 856
rect 213846 734 214322 856
rect 214490 734 214966 856
rect 215134 734 215610 856
rect 215778 734 216254 856
rect 216422 734 216898 856
rect 217066 734 217542 856
rect 217710 734 218186 856
rect 218354 734 218830 856
rect 218998 734 219474 856
rect 219642 734 220118 856
rect 220286 734 220762 856
rect 220930 734 221406 856
rect 221574 734 222050 856
rect 222218 734 222694 856
rect 222862 734 223338 856
rect 223506 734 223982 856
rect 224150 734 224626 856
rect 224794 734 225270 856
rect 225438 734 225914 856
rect 226082 734 226558 856
rect 226726 734 227202 856
rect 227370 734 227846 856
rect 228014 734 228490 856
rect 228658 734 229134 856
rect 229302 734 229778 856
rect 229946 734 230422 856
rect 230590 734 231066 856
rect 231234 734 231710 856
rect 231878 734 232354 856
rect 232522 734 232998 856
rect 233166 734 233642 856
rect 233810 734 234286 856
rect 234454 734 234930 856
rect 235098 734 235574 856
rect 235742 734 236218 856
rect 236386 734 236862 856
rect 237030 734 237506 856
rect 237674 734 238150 856
rect 238318 734 238794 856
rect 238962 734 239438 856
rect 239606 734 240082 856
rect 240250 734 240726 856
rect 240894 734 241370 856
rect 241538 734 242014 856
rect 242182 734 242658 856
rect 242826 734 243302 856
rect 243470 734 243946 856
rect 244114 734 244590 856
rect 244758 734 245234 856
rect 245402 734 245878 856
rect 246046 734 246522 856
rect 246690 734 247166 856
rect 247334 734 247810 856
rect 247978 734 248454 856
rect 248622 734 249098 856
rect 249266 734 249742 856
rect 249910 734 250386 856
rect 250554 734 251030 856
rect 251198 734 251674 856
rect 251842 734 252318 856
rect 252486 734 252962 856
rect 253130 734 253606 856
rect 253774 734 254250 856
rect 254418 734 254894 856
rect 255062 734 255538 856
rect 255706 734 256182 856
rect 256350 734 256826 856
rect 256994 734 257470 856
rect 257638 734 258114 856
rect 258282 734 258758 856
rect 258926 734 259402 856
rect 259570 734 260046 856
rect 260214 734 260690 856
rect 260858 734 261334 856
rect 261502 734 261978 856
rect 262146 734 262622 856
rect 262790 734 263266 856
rect 263434 734 263910 856
rect 264078 734 264554 856
rect 264722 734 265198 856
rect 265366 734 265842 856
rect 266010 734 266486 856
rect 266654 734 267130 856
rect 267298 734 267774 856
rect 267942 734 268418 856
rect 268586 734 269062 856
rect 269230 734 269706 856
rect 269874 734 270350 856
rect 270518 734 270994 856
rect 271162 734 271638 856
rect 271806 734 272282 856
rect 272450 734 272926 856
rect 273094 734 273570 856
rect 273738 734 274214 856
rect 274382 734 274858 856
rect 275026 734 275502 856
rect 275670 734 276146 856
rect 276314 734 276790 856
rect 276958 734 277434 856
rect 277602 734 278078 856
rect 278246 734 278722 856
rect 278890 734 279366 856
rect 279534 734 280010 856
rect 280178 734 280654 856
rect 280822 734 281298 856
rect 281466 734 281942 856
rect 282110 734 282586 856
rect 282754 734 283230 856
rect 283398 734 283874 856
rect 284042 734 284518 856
rect 284686 734 285162 856
rect 285330 734 285806 856
rect 285974 734 286450 856
rect 286618 734 287094 856
rect 287262 734 287738 856
rect 287906 734 288382 856
rect 288550 734 289026 856
rect 289194 734 289670 856
rect 289838 734 290314 856
rect 290482 734 290958 856
rect 291126 734 291602 856
rect 291770 734 292246 856
rect 292414 734 292890 856
rect 293058 734 293534 856
rect 293702 734 294178 856
rect 294346 734 294822 856
rect 294990 734 295466 856
rect 295634 734 296110 856
rect 296278 734 296754 856
rect 296922 734 297398 856
rect 297566 734 298042 856
rect 298210 734 298686 856
rect 298854 734 299330 856
rect 299498 734 299974 856
rect 300142 734 300618 856
rect 300786 734 301262 856
rect 301430 734 301906 856
rect 302074 734 302550 856
rect 302718 734 303194 856
rect 303362 734 303838 856
rect 304006 734 304482 856
rect 304650 734 305126 856
rect 305294 734 305770 856
rect 305938 734 306414 856
rect 306582 734 307058 856
rect 307226 734 307702 856
rect 307870 734 308346 856
rect 308514 734 308990 856
rect 309158 734 309634 856
rect 309802 734 310278 856
rect 310446 734 310922 856
rect 311090 734 311566 856
rect 311734 734 312210 856
rect 312378 734 312854 856
rect 313022 734 313498 856
rect 313666 734 314142 856
rect 314310 734 314786 856
rect 314954 734 315430 856
rect 315598 734 316074 856
rect 316242 734 316718 856
rect 316886 734 317362 856
rect 317530 734 318006 856
rect 318174 734 318650 856
<< metal3 >>
rect 319200 315528 320000 315648
rect 0 314848 800 314968
rect 319200 309544 320000 309664
rect 0 309000 800 309120
rect 319200 303560 320000 303680
rect 0 303152 800 303272
rect 319200 297576 320000 297696
rect 0 297304 800 297424
rect 0 291456 800 291576
rect 319200 291592 320000 291712
rect 0 285608 800 285728
rect 319200 285608 320000 285728
rect 0 279760 800 279880
rect 319200 279624 320000 279744
rect 0 273912 800 274032
rect 319200 273640 320000 273760
rect 0 268064 800 268184
rect 319200 267656 320000 267776
rect 0 262216 800 262336
rect 319200 261672 320000 261792
rect 0 256368 800 256488
rect 319200 255688 320000 255808
rect 0 250520 800 250640
rect 319200 249704 320000 249824
rect 0 244672 800 244792
rect 319200 243720 320000 243840
rect 0 238824 800 238944
rect 319200 237736 320000 237856
rect 0 232976 800 233096
rect 319200 231752 320000 231872
rect 0 227128 800 227248
rect 319200 225768 320000 225888
rect 0 221280 800 221400
rect 319200 219784 320000 219904
rect 0 215432 800 215552
rect 319200 213800 320000 213920
rect 0 209584 800 209704
rect 319200 207816 320000 207936
rect 0 203736 800 203856
rect 319200 201832 320000 201952
rect 0 197888 800 198008
rect 319200 195848 320000 195968
rect 0 192040 800 192160
rect 319200 189864 320000 189984
rect 0 186192 800 186312
rect 319200 183880 320000 184000
rect 0 180344 800 180464
rect 319200 177896 320000 178016
rect 0 174496 800 174616
rect 319200 171912 320000 172032
rect 0 168648 800 168768
rect 319200 165928 320000 166048
rect 0 162800 800 162920
rect 319200 159944 320000 160064
rect 0 156952 800 157072
rect 319200 153960 320000 154080
rect 0 151104 800 151224
rect 319200 147976 320000 148096
rect 0 145256 800 145376
rect 319200 141992 320000 142112
rect 0 139408 800 139528
rect 319200 136008 320000 136128
rect 0 133560 800 133680
rect 319200 130024 320000 130144
rect 0 127712 800 127832
rect 319200 124040 320000 124160
rect 0 121864 800 121984
rect 319200 118056 320000 118176
rect 0 116016 800 116136
rect 319200 112072 320000 112192
rect 0 110168 800 110288
rect 319200 106088 320000 106208
rect 0 104320 800 104440
rect 319200 100104 320000 100224
rect 0 98472 800 98592
rect 319200 94120 320000 94240
rect 0 92624 800 92744
rect 319200 88136 320000 88256
rect 0 86776 800 86896
rect 319200 82152 320000 82272
rect 0 80928 800 81048
rect 319200 76168 320000 76288
rect 0 75080 800 75200
rect 319200 70184 320000 70304
rect 0 69232 800 69352
rect 319200 64200 320000 64320
rect 0 63384 800 63504
rect 319200 58216 320000 58336
rect 0 57536 800 57656
rect 319200 52232 320000 52352
rect 0 51688 800 51808
rect 319200 46248 320000 46368
rect 0 45840 800 45960
rect 319200 40264 320000 40384
rect 0 39992 800 40112
rect 0 34144 800 34264
rect 319200 34280 320000 34400
rect 0 28296 800 28416
rect 319200 28296 320000 28416
rect 0 22448 800 22568
rect 319200 22312 320000 22432
rect 0 16600 800 16720
rect 319200 16328 320000 16448
rect 0 10752 800 10872
rect 319200 10344 320000 10464
rect 0 4904 800 5024
rect 319200 4360 320000 4480
<< obsm3 >>
rect 800 315728 319200 317729
rect 800 315448 319120 315728
rect 800 315048 319200 315448
rect 880 314768 319200 315048
rect 800 309744 319200 314768
rect 800 309464 319120 309744
rect 800 309200 319200 309464
rect 880 308920 319200 309200
rect 800 303760 319200 308920
rect 800 303480 319120 303760
rect 800 303352 319200 303480
rect 880 303072 319200 303352
rect 800 297776 319200 303072
rect 800 297504 319120 297776
rect 880 297496 319120 297504
rect 880 297224 319200 297496
rect 800 291792 319200 297224
rect 800 291656 319120 291792
rect 880 291512 319120 291656
rect 880 291376 319200 291512
rect 800 285808 319200 291376
rect 880 285528 319120 285808
rect 800 279960 319200 285528
rect 880 279824 319200 279960
rect 880 279680 319120 279824
rect 800 279544 319120 279680
rect 800 274112 319200 279544
rect 880 273840 319200 274112
rect 880 273832 319120 273840
rect 800 273560 319120 273832
rect 800 268264 319200 273560
rect 880 267984 319200 268264
rect 800 267856 319200 267984
rect 800 267576 319120 267856
rect 800 262416 319200 267576
rect 880 262136 319200 262416
rect 800 261872 319200 262136
rect 800 261592 319120 261872
rect 800 256568 319200 261592
rect 880 256288 319200 256568
rect 800 255888 319200 256288
rect 800 255608 319120 255888
rect 800 250720 319200 255608
rect 880 250440 319200 250720
rect 800 249904 319200 250440
rect 800 249624 319120 249904
rect 800 244872 319200 249624
rect 880 244592 319200 244872
rect 800 243920 319200 244592
rect 800 243640 319120 243920
rect 800 239024 319200 243640
rect 880 238744 319200 239024
rect 800 237936 319200 238744
rect 800 237656 319120 237936
rect 800 233176 319200 237656
rect 880 232896 319200 233176
rect 800 231952 319200 232896
rect 800 231672 319120 231952
rect 800 227328 319200 231672
rect 880 227048 319200 227328
rect 800 225968 319200 227048
rect 800 225688 319120 225968
rect 800 221480 319200 225688
rect 880 221200 319200 221480
rect 800 219984 319200 221200
rect 800 219704 319120 219984
rect 800 215632 319200 219704
rect 880 215352 319200 215632
rect 800 214000 319200 215352
rect 800 213720 319120 214000
rect 800 209784 319200 213720
rect 880 209504 319200 209784
rect 800 208016 319200 209504
rect 800 207736 319120 208016
rect 800 203936 319200 207736
rect 880 203656 319200 203936
rect 800 202032 319200 203656
rect 800 201752 319120 202032
rect 800 198088 319200 201752
rect 880 197808 319200 198088
rect 800 196048 319200 197808
rect 800 195768 319120 196048
rect 800 192240 319200 195768
rect 880 191960 319200 192240
rect 800 190064 319200 191960
rect 800 189784 319120 190064
rect 800 186392 319200 189784
rect 880 186112 319200 186392
rect 800 184080 319200 186112
rect 800 183800 319120 184080
rect 800 180544 319200 183800
rect 880 180264 319200 180544
rect 800 178096 319200 180264
rect 800 177816 319120 178096
rect 800 174696 319200 177816
rect 880 174416 319200 174696
rect 800 172112 319200 174416
rect 800 171832 319120 172112
rect 800 168848 319200 171832
rect 880 168568 319200 168848
rect 800 166128 319200 168568
rect 800 165848 319120 166128
rect 800 163000 319200 165848
rect 880 162720 319200 163000
rect 800 160144 319200 162720
rect 800 159864 319120 160144
rect 800 157152 319200 159864
rect 880 156872 319200 157152
rect 800 154160 319200 156872
rect 800 153880 319120 154160
rect 800 151304 319200 153880
rect 880 151024 319200 151304
rect 800 148176 319200 151024
rect 800 147896 319120 148176
rect 800 145456 319200 147896
rect 880 145176 319200 145456
rect 800 142192 319200 145176
rect 800 141912 319120 142192
rect 800 139608 319200 141912
rect 880 139328 319200 139608
rect 800 136208 319200 139328
rect 800 135928 319120 136208
rect 800 133760 319200 135928
rect 880 133480 319200 133760
rect 800 130224 319200 133480
rect 800 129944 319120 130224
rect 800 127912 319200 129944
rect 880 127632 319200 127912
rect 800 124240 319200 127632
rect 800 123960 319120 124240
rect 800 122064 319200 123960
rect 880 121784 319200 122064
rect 800 118256 319200 121784
rect 800 117976 319120 118256
rect 800 116216 319200 117976
rect 880 115936 319200 116216
rect 800 112272 319200 115936
rect 800 111992 319120 112272
rect 800 110368 319200 111992
rect 880 110088 319200 110368
rect 800 106288 319200 110088
rect 800 106008 319120 106288
rect 800 104520 319200 106008
rect 880 104240 319200 104520
rect 800 100304 319200 104240
rect 800 100024 319120 100304
rect 800 98672 319200 100024
rect 880 98392 319200 98672
rect 800 94320 319200 98392
rect 800 94040 319120 94320
rect 800 92824 319200 94040
rect 880 92544 319200 92824
rect 800 88336 319200 92544
rect 800 88056 319120 88336
rect 800 86976 319200 88056
rect 880 86696 319200 86976
rect 800 82352 319200 86696
rect 800 82072 319120 82352
rect 800 81128 319200 82072
rect 880 80848 319200 81128
rect 800 76368 319200 80848
rect 800 76088 319120 76368
rect 800 75280 319200 76088
rect 880 75000 319200 75280
rect 800 70384 319200 75000
rect 800 70104 319120 70384
rect 800 69432 319200 70104
rect 880 69152 319200 69432
rect 800 64400 319200 69152
rect 800 64120 319120 64400
rect 800 63584 319200 64120
rect 880 63304 319200 63584
rect 800 58416 319200 63304
rect 800 58136 319120 58416
rect 800 57736 319200 58136
rect 880 57456 319200 57736
rect 800 52432 319200 57456
rect 800 52152 319120 52432
rect 800 51888 319200 52152
rect 880 51608 319200 51888
rect 800 46448 319200 51608
rect 800 46168 319120 46448
rect 800 46040 319200 46168
rect 880 45760 319200 46040
rect 800 40464 319200 45760
rect 800 40192 319120 40464
rect 880 40184 319120 40192
rect 880 39912 319200 40184
rect 800 34480 319200 39912
rect 800 34344 319120 34480
rect 880 34200 319120 34344
rect 880 34064 319200 34200
rect 800 28496 319200 34064
rect 880 28216 319120 28496
rect 800 22648 319200 28216
rect 880 22512 319200 22648
rect 880 22368 319120 22512
rect 800 22232 319120 22368
rect 800 16800 319200 22232
rect 880 16528 319200 16800
rect 880 16520 319120 16528
rect 800 16248 319120 16520
rect 800 10952 319200 16248
rect 880 10672 319200 10952
rect 800 10544 319200 10672
rect 800 10264 319120 10544
rect 800 5104 319200 10264
rect 880 4824 319200 5104
rect 800 4560 319200 4824
rect 800 4280 319120 4560
rect 800 2143 319200 4280
<< metal4 >>
rect 4208 2128 4528 317744
rect 4868 2128 5188 317744
rect 34928 2128 35248 317744
rect 35588 2128 35908 317744
rect 65648 2128 65968 317744
rect 66308 2128 66628 317744
rect 96368 2128 96688 317744
rect 97028 2128 97348 317744
rect 127088 2128 127408 317744
rect 127748 2128 128068 317744
rect 157808 2128 158128 317744
rect 158468 2128 158788 317744
rect 188528 2128 188848 317744
rect 189188 2128 189508 317744
rect 219248 2128 219568 317744
rect 219908 2128 220228 317744
rect 249968 2128 250288 317744
rect 250628 2128 250948 317744
rect 280688 2128 281008 317744
rect 281348 2128 281668 317744
rect 311408 2128 311728 317744
rect 312068 2128 312388 317744
<< obsm4 >>
rect 259499 215051 280608 317525
rect 281088 215051 281268 317525
rect 281748 215051 311328 317525
rect 311808 215051 311988 317525
rect 312468 215051 314213 317525
<< metal5 >>
rect 1056 312366 318920 312686
rect 1056 311706 318920 312026
rect 1056 281730 318920 282050
rect 1056 281070 318920 281390
rect 1056 251094 318920 251414
rect 1056 250434 318920 250754
rect 1056 220458 318920 220778
rect 1056 219798 318920 220118
rect 1056 189822 318920 190142
rect 1056 189162 318920 189482
rect 1056 159186 318920 159506
rect 1056 158526 318920 158846
rect 1056 128550 318920 128870
rect 1056 127890 318920 128210
rect 1056 97914 318920 98234
rect 1056 97254 318920 97574
rect 1056 67278 318920 67598
rect 1056 66618 318920 66938
rect 1056 36642 318920 36962
rect 1056 35982 318920 36302
rect 1056 6006 318920 6326
rect 1056 5346 318920 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127748 2128 128068 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 158468 2128 158788 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 189188 2128 189508 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 219908 2128 220228 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 250628 2128 250948 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 281348 2128 281668 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 312068 2128 312388 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 318920 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 318920 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 318920 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 318920 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 128550 318920 128870 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 159186 318920 159506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 189822 318920 190142 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 220458 318920 220778 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 251094 318920 251414 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 281730 318920 282050 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 312366 318920 312686 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 318920 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 318920 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 318920 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 318920 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 318920 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 158526 318920 158846 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 189162 318920 189482 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 219798 318920 220118 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 250434 318920 250754 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 281070 318920 281390 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 311706 318920 312026 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 319200 130024 320000 130144 6 analog_io[0]
port 3 nsew signal bidirectional
rlabel metal2 s 243818 319200 243874 320000 6 analog_io[10]
port 4 nsew signal bidirectional
rlabel metal2 s 208490 319200 208546 320000 6 analog_io[11]
port 5 nsew signal bidirectional
rlabel metal2 s 173162 319200 173218 320000 6 analog_io[12]
port 6 nsew signal bidirectional
rlabel metal2 s 137834 319200 137890 320000 6 analog_io[13]
port 7 nsew signal bidirectional
rlabel metal2 s 102506 319200 102562 320000 6 analog_io[14]
port 8 nsew signal bidirectional
rlabel metal2 s 67178 319200 67234 320000 6 analog_io[15]
port 9 nsew signal bidirectional
rlabel metal2 s 31850 319200 31906 320000 6 analog_io[16]
port 10 nsew signal bidirectional
rlabel metal3 s 0 314848 800 314968 6 analog_io[17]
port 11 nsew signal bidirectional
rlabel metal3 s 0 291456 800 291576 6 analog_io[18]
port 12 nsew signal bidirectional
rlabel metal3 s 0 268064 800 268184 6 analog_io[19]
port 13 nsew signal bidirectional
rlabel metal3 s 319200 153960 320000 154080 6 analog_io[1]
port 14 nsew signal bidirectional
rlabel metal3 s 0 244672 800 244792 6 analog_io[20]
port 15 nsew signal bidirectional
rlabel metal3 s 0 221280 800 221400 6 analog_io[21]
port 16 nsew signal bidirectional
rlabel metal3 s 0 197888 800 198008 6 analog_io[22]
port 17 nsew signal bidirectional
rlabel metal3 s 0 174496 800 174616 6 analog_io[23]
port 18 nsew signal bidirectional
rlabel metal3 s 0 151104 800 151224 6 analog_io[24]
port 19 nsew signal bidirectional
rlabel metal3 s 0 127712 800 127832 6 analog_io[25]
port 20 nsew signal bidirectional
rlabel metal3 s 0 104320 800 104440 6 analog_io[26]
port 21 nsew signal bidirectional
rlabel metal3 s 0 80928 800 81048 6 analog_io[27]
port 22 nsew signal bidirectional
rlabel metal3 s 0 57536 800 57656 6 analog_io[28]
port 23 nsew signal bidirectional
rlabel metal3 s 319200 177896 320000 178016 6 analog_io[2]
port 24 nsew signal bidirectional
rlabel metal3 s 319200 201832 320000 201952 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 319200 225768 320000 225888 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 319200 249704 320000 249824 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 319200 273640 320000 273760 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 319200 297576 320000 297696 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 314474 319200 314530 320000 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 279146 319200 279202 320000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal3 s 319200 4360 320000 4480 6 io_in[0]
port 32 nsew signal input
rlabel metal3 s 319200 207816 320000 207936 6 io_in[10]
port 33 nsew signal input
rlabel metal3 s 319200 231752 320000 231872 6 io_in[11]
port 34 nsew signal input
rlabel metal3 s 319200 255688 320000 255808 6 io_in[12]
port 35 nsew signal input
rlabel metal3 s 319200 279624 320000 279744 6 io_in[13]
port 36 nsew signal input
rlabel metal3 s 319200 303560 320000 303680 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 305642 319200 305698 320000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 270314 319200 270370 320000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 234986 319200 235042 320000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 199658 319200 199714 320000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 164330 319200 164386 320000 6 io_in[19]
port 42 nsew signal input
rlabel metal3 s 319200 22312 320000 22432 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 129002 319200 129058 320000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 93674 319200 93730 320000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 58346 319200 58402 320000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 23018 319200 23074 320000 6 io_in[23]
port 47 nsew signal input
rlabel metal3 s 0 309000 800 309120 6 io_in[24]
port 48 nsew signal input
rlabel metal3 s 0 285608 800 285728 6 io_in[25]
port 49 nsew signal input
rlabel metal3 s 0 262216 800 262336 6 io_in[26]
port 50 nsew signal input
rlabel metal3 s 0 238824 800 238944 6 io_in[27]
port 51 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 io_in[28]
port 52 nsew signal input
rlabel metal3 s 0 192040 800 192160 6 io_in[29]
port 53 nsew signal input
rlabel metal3 s 319200 40264 320000 40384 6 io_in[2]
port 54 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 io_in[30]
port 55 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 io_in[31]
port 56 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 io_in[32]
port 57 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 io_in[33]
port 58 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 io_in[34]
port 59 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_in[35]
port 60 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 io_in[36]
port 61 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[37]
port 62 nsew signal input
rlabel metal3 s 319200 58216 320000 58336 6 io_in[3]
port 63 nsew signal input
rlabel metal3 s 319200 76168 320000 76288 6 io_in[4]
port 64 nsew signal input
rlabel metal3 s 319200 94120 320000 94240 6 io_in[5]
port 65 nsew signal input
rlabel metal3 s 319200 112072 320000 112192 6 io_in[6]
port 66 nsew signal input
rlabel metal3 s 319200 136008 320000 136128 6 io_in[7]
port 67 nsew signal input
rlabel metal3 s 319200 159944 320000 160064 6 io_in[8]
port 68 nsew signal input
rlabel metal3 s 319200 183880 320000 184000 6 io_in[9]
port 69 nsew signal input
rlabel metal3 s 319200 16328 320000 16448 6 io_oeb[0]
port 70 nsew signal output
rlabel metal3 s 319200 219784 320000 219904 6 io_oeb[10]
port 71 nsew signal output
rlabel metal3 s 319200 243720 320000 243840 6 io_oeb[11]
port 72 nsew signal output
rlabel metal3 s 319200 267656 320000 267776 6 io_oeb[12]
port 73 nsew signal output
rlabel metal3 s 319200 291592 320000 291712 6 io_oeb[13]
port 74 nsew signal output
rlabel metal3 s 319200 315528 320000 315648 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 287978 319200 288034 320000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 252650 319200 252706 320000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 217322 319200 217378 320000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 181994 319200 182050 320000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 146666 319200 146722 320000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal3 s 319200 34280 320000 34400 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 111338 319200 111394 320000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 76010 319200 76066 320000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 40682 319200 40738 320000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 5354 319200 5410 320000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal3 s 0 297304 800 297424 6 io_oeb[24]
port 86 nsew signal output
rlabel metal3 s 0 273912 800 274032 6 io_oeb[25]
port 87 nsew signal output
rlabel metal3 s 0 250520 800 250640 6 io_oeb[26]
port 88 nsew signal output
rlabel metal3 s 0 227128 800 227248 6 io_oeb[27]
port 89 nsew signal output
rlabel metal3 s 0 203736 800 203856 6 io_oeb[28]
port 90 nsew signal output
rlabel metal3 s 0 180344 800 180464 6 io_oeb[29]
port 91 nsew signal output
rlabel metal3 s 319200 52232 320000 52352 6 io_oeb[2]
port 92 nsew signal output
rlabel metal3 s 0 156952 800 157072 6 io_oeb[30]
port 93 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 io_oeb[31]
port 94 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 io_oeb[32]
port 95 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 io_oeb[33]
port 96 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 io_oeb[34]
port 97 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 io_oeb[35]
port 98 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 io_oeb[36]
port 99 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 io_oeb[37]
port 100 nsew signal output
rlabel metal3 s 319200 70184 320000 70304 6 io_oeb[3]
port 101 nsew signal output
rlabel metal3 s 319200 88136 320000 88256 6 io_oeb[4]
port 102 nsew signal output
rlabel metal3 s 319200 106088 320000 106208 6 io_oeb[5]
port 103 nsew signal output
rlabel metal3 s 319200 124040 320000 124160 6 io_oeb[6]
port 104 nsew signal output
rlabel metal3 s 319200 147976 320000 148096 6 io_oeb[7]
port 105 nsew signal output
rlabel metal3 s 319200 171912 320000 172032 6 io_oeb[8]
port 106 nsew signal output
rlabel metal3 s 319200 195848 320000 195968 6 io_oeb[9]
port 107 nsew signal output
rlabel metal3 s 319200 10344 320000 10464 6 io_out[0]
port 108 nsew signal output
rlabel metal3 s 319200 213800 320000 213920 6 io_out[10]
port 109 nsew signal output
rlabel metal3 s 319200 237736 320000 237856 6 io_out[11]
port 110 nsew signal output
rlabel metal3 s 319200 261672 320000 261792 6 io_out[12]
port 111 nsew signal output
rlabel metal3 s 319200 285608 320000 285728 6 io_out[13]
port 112 nsew signal output
rlabel metal3 s 319200 309544 320000 309664 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 296810 319200 296866 320000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 261482 319200 261538 320000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 226154 319200 226210 320000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 190826 319200 190882 320000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 155498 319200 155554 320000 6 io_out[19]
port 118 nsew signal output
rlabel metal3 s 319200 28296 320000 28416 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 120170 319200 120226 320000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 84842 319200 84898 320000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 49514 319200 49570 320000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 14186 319200 14242 320000 6 io_out[23]
port 123 nsew signal output
rlabel metal3 s 0 303152 800 303272 6 io_out[24]
port 124 nsew signal output
rlabel metal3 s 0 279760 800 279880 6 io_out[25]
port 125 nsew signal output
rlabel metal3 s 0 256368 800 256488 6 io_out[26]
port 126 nsew signal output
rlabel metal3 s 0 232976 800 233096 6 io_out[27]
port 127 nsew signal output
rlabel metal3 s 0 209584 800 209704 6 io_out[28]
port 128 nsew signal output
rlabel metal3 s 0 186192 800 186312 6 io_out[29]
port 129 nsew signal output
rlabel metal3 s 319200 46248 320000 46368 6 io_out[2]
port 130 nsew signal output
rlabel metal3 s 0 162800 800 162920 6 io_out[30]
port 131 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 io_out[31]
port 132 nsew signal output
rlabel metal3 s 0 116016 800 116136 6 io_out[32]
port 133 nsew signal output
rlabel metal3 s 0 92624 800 92744 6 io_out[33]
port 134 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 io_out[34]
port 135 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_out[35]
port 136 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 io_out[36]
port 137 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 io_out[37]
port 138 nsew signal output
rlabel metal3 s 319200 64200 320000 64320 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 319200 82152 320000 82272 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 319200 100104 320000 100224 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 319200 118056 320000 118176 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 319200 141992 320000 142112 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 319200 165928 320000 166048 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 319200 189864 320000 189984 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 276202 0 276258 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 280066 0 280122 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 283930 0 283986 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 285862 0 285918 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 287794 0 287850 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 291658 0 291714 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 293590 0 293646 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 295522 0 295578 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 297454 0 297510 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 301318 0 301374 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 303250 0 303306 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 305182 0 305238 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 307114 0 307170 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 309046 0 309102 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 310978 0 311034 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 312910 0 312966 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 314842 0 314898 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 193126 0 193182 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 220174 0 220230 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 239494 0 239550 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 241426 0 241482 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 256882 0 256938 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 263322 0 263378 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 265254 0 265310 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 267186 0 267242 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 269118 0 269174 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 271050 0 271106 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 272982 0 273038 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 274914 0 274970 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 276846 0 276902 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 280710 0 280766 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 282642 0 282698 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 284574 0 284630 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 286506 0 286562 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 288438 0 288494 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 290370 0 290426 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 292302 0 292358 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 294234 0 294290 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 296166 0 296222 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 298098 0 298154 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 300030 0 300086 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 301962 0 302018 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 303894 0 303950 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 305826 0 305882 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 307758 0 307814 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 309690 0 309746 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 311622 0 311678 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 315486 0 315542 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 158994 0 159050 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 168654 0 168710 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 193770 0 193826 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 197634 0 197690 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 199566 0 199622 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 203430 0 203486 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 205362 0 205418 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 207294 0 207350 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 213090 0 213146 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 216954 0 217010 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 220818 0 220874 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 224682 0 224738 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 226614 0 226670 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 228546 0 228602 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 232410 0 232466 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 238206 0 238262 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 242070 0 242126 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 247866 0 247922 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 249798 0 249854 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 253662 0 253718 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 255594 0 255650 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 257526 0 257582 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 259458 0 259514 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 261390 0 261446 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_oenb[0]
port 402 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_oenb[100]
port 403 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_oenb[101]
port 404 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_oenb[102]
port 405 nsew signal input
rlabel metal2 s 269762 0 269818 800 6 la_oenb[103]
port 406 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_oenb[104]
port 407 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_oenb[105]
port 408 nsew signal input
rlabel metal2 s 275558 0 275614 800 6 la_oenb[106]
port 409 nsew signal input
rlabel metal2 s 277490 0 277546 800 6 la_oenb[107]
port 410 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oenb[108]
port 411 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_oenb[109]
port 412 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[10]
port 413 nsew signal input
rlabel metal2 s 283286 0 283342 800 6 la_oenb[110]
port 414 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_oenb[111]
port 415 nsew signal input
rlabel metal2 s 287150 0 287206 800 6 la_oenb[112]
port 416 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_oenb[113]
port 417 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_oenb[114]
port 418 nsew signal input
rlabel metal2 s 292946 0 293002 800 6 la_oenb[115]
port 419 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[116]
port 420 nsew signal input
rlabel metal2 s 296810 0 296866 800 6 la_oenb[117]
port 421 nsew signal input
rlabel metal2 s 298742 0 298798 800 6 la_oenb[118]
port 422 nsew signal input
rlabel metal2 s 300674 0 300730 800 6 la_oenb[119]
port 423 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[11]
port 424 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_oenb[120]
port 425 nsew signal input
rlabel metal2 s 304538 0 304594 800 6 la_oenb[121]
port 426 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_oenb[122]
port 427 nsew signal input
rlabel metal2 s 308402 0 308458 800 6 la_oenb[123]
port 428 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_oenb[124]
port 429 nsew signal input
rlabel metal2 s 312266 0 312322 800 6 la_oenb[125]
port 430 nsew signal input
rlabel metal2 s 314198 0 314254 800 6 la_oenb[126]
port 431 nsew signal input
rlabel metal2 s 316130 0 316186 800 6 la_oenb[127]
port 432 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[12]
port 433 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[13]
port 434 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[14]
port 435 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[15]
port 436 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[16]
port 437 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[17]
port 438 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_oenb[18]
port 439 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[19]
port 440 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[1]
port 441 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[20]
port 442 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[21]
port 443 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[22]
port 444 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_oenb[23]
port 445 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[24]
port 446 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[25]
port 447 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_oenb[26]
port 448 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[27]
port 449 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[28]
port 450 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[29]
port 451 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[2]
port 452 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[30]
port 453 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[31]
port 454 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[32]
port 455 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[33]
port 456 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[34]
port 457 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[35]
port 458 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[36]
port 459 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[37]
port 460 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[38]
port 461 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[39]
port 462 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[3]
port 463 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[40]
port 464 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[41]
port 465 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[42]
port 466 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[43]
port 467 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_oenb[44]
port 468 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_oenb[45]
port 469 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[46]
port 470 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[47]
port 471 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_oenb[48]
port 472 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oenb[49]
port 473 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[4]
port 474 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[50]
port 475 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_oenb[51]
port 476 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[52]
port 477 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[53]
port 478 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_oenb[54]
port 479 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_oenb[55]
port 480 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[56]
port 481 nsew signal input
rlabel metal2 s 180890 0 180946 800 6 la_oenb[57]
port 482 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_oenb[58]
port 483 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_oenb[59]
port 484 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[5]
port 485 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_oenb[60]
port 486 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oenb[61]
port 487 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_oenb[62]
port 488 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_oenb[63]
port 489 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oenb[64]
port 490 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oenb[65]
port 491 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_oenb[66]
port 492 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_oenb[67]
port 493 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_oenb[68]
port 494 nsew signal input
rlabel metal2 s 204074 0 204130 800 6 la_oenb[69]
port 495 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[6]
port 496 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_oenb[70]
port 497 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_oenb[71]
port 498 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[72]
port 499 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_oenb[73]
port 500 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_oenb[74]
port 501 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_oenb[75]
port 502 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_oenb[76]
port 503 nsew signal input
rlabel metal2 s 219530 0 219586 800 6 la_oenb[77]
port 504 nsew signal input
rlabel metal2 s 221462 0 221518 800 6 la_oenb[78]
port 505 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_oenb[79]
port 506 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[7]
port 507 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_oenb[80]
port 508 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_oenb[81]
port 509 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 la_oenb[82]
port 510 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oenb[83]
port 511 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_oenb[84]
port 512 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_oenb[85]
port 513 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[86]
port 514 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oenb[87]
port 515 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_oenb[88]
port 516 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_oenb[89]
port 517 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[8]
port 518 nsew signal input
rlabel metal2 s 244646 0 244702 800 6 la_oenb[90]
port 519 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_oenb[91]
port 520 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_oenb[92]
port 521 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_oenb[93]
port 522 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_oenb[94]
port 523 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_oenb[95]
port 524 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oenb[96]
port 525 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oenb[97]
port 526 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oenb[98]
port 527 nsew signal input
rlabel metal2 s 262034 0 262090 800 6 la_oenb[99]
port 528 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[9]
port 529 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 317418 0 317474 800 6 user_irq[0]
port 531 nsew signal output
rlabel metal2 s 318062 0 318118 800 6 user_irq[1]
port 532 nsew signal output
rlabel metal2 s 318706 0 318762 800 6 user_irq[2]
port 533 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 39130774
string GDS_FILE /openlane/designs/pipeline_mul_tapeout/runs/RUN_2023.11.25_16.31.35/results/signoff/user_project_wrapper.magic.gds
string GDS_START 892612
<< end >>

